module MIYAJIRO_CPU(
    input reset_n,
    input clk
);

endmodule
